// Register with enabled and async reset
module floper #(
    parameter int Width = 1,
    parameter logic[Width-1:0] ResetValue = '0
)(
    input logic clk, reset_n, en,
    input logic[Width-1:0] d,
    output logic[Width-1:0] q
);
    always_ff @(posedge clk or negedge reset_n) begin
        if (~reset_n) q <= ResetValue;
        else if (en) q <= d;
    end
endmodule
